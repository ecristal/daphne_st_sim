module st40_top_wrapper(
    input wire reset_aclk,
    input wire reset_fclk,
    input wire [7:0] adhoc,
    input wire [13:0] st_config,
    input wire [4:0] signal_delay,
    input wire [41:0] threshold_xc,
    input wire [7:0] ti_trigger,
    input wire ti_trigger_stbr,
    input wire reset_st_counters,
    input wire [3:0] slot_id,
    input wire [9:0] crate_id,
    input wire [5:0] detector_id,
    input wire [5:0] version_id,
    input wire [39:0] enable,
    input wire [39:0] afe_comp_enable,
    input wire [39:0] invert_enable,
    input wire [5:0] st_40_signals_enable_reg,
    output wire st_40_selftrigger_4_spybuffer,
    input wire [1:0] filter_output_selector,
    input wire aclk,
    input wire [63:0] timestamp,
    input wire [13:0] afe_dat_0_0,
    input wire [13:0] afe_dat_0_1,
    input wire [13:0] afe_dat_0_2,
    input wire [13:0] afe_dat_0_3,
    input wire [13:0] afe_dat_0_4,
    input wire [13:0] afe_dat_0_5,
    input wire [13:0] afe_dat_0_6,
    input wire [13:0] afe_dat_0_7,
    input wire [13:0] afe_dat_0_8,
    input wire [13:0] afe_dat_1_0,
    input wire [13:0] afe_dat_1_1,
    input wire [13:0] afe_dat_1_2,
    input wire [13:0] afe_dat_1_3,
    input wire [13:0] afe_dat_1_4,
    input wire [13:0] afe_dat_1_5,
    input wire [13:0] afe_dat_1_6,
    input wire [13:0] afe_dat_1_7,
    input wire [13:0] afe_dat_1_8,
    input wire [13:0] afe_dat_2_0,
    input wire [13:0] afe_dat_2_1,
    input wire [13:0] afe_dat_2_2,
    input wire [13:0] afe_dat_2_3,
    input wire [13:0] afe_dat_2_4,
    input wire [13:0] afe_dat_2_5,
    input wire [13:0] afe_dat_2_6,
    input wire [13:0] afe_dat_2_7,
    input wire [13:0] afe_dat_2_8,
    input wire [13:0] afe_dat_3_0,
    input wire [13:0] afe_dat_3_1,
    input wire [13:0] afe_dat_3_2,
    input wire [13:0] afe_dat_3_3,
    input wire [13:0] afe_dat_3_4,
    input wire [13:0] afe_dat_3_5,
    input wire [13:0] afe_dat_3_6,
    input wire [13:0] afe_dat_3_7,
    input wire [13:0] afe_dat_3_8,
    input wire [13:0] afe_dat_4_0,
    input wire [13:0] afe_dat_4_1,
    input wire [13:0] afe_dat_4_2,
    input wire [13:0] afe_dat_4_3,
    input wire [13:0] afe_dat_4_4,
    input wire [13:0] afe_dat_4_5,
    input wire [13:0] afe_dat_4_6,
    input wire [13:0] afe_dat_4_7,
    input wire [13:0] afe_dat_4_8,
    output wire [13:0] afe_dat_0_0_filtered,
    output wire [13:0] afe_dat_0_1_filtered,
    output wire [13:0] afe_dat_0_2_filtered,
    output wire [13:0] afe_dat_0_3_filtered,
    output wire [13:0] afe_dat_0_4_filtered,
    output wire [13:0] afe_dat_0_5_filtered,
    output wire [13:0] afe_dat_0_6_filtered,
    output wire [13:0] afe_dat_0_7_filtered,
    output wire [13:0] afe_dat_0_8_filtered,
    output wire [13:0] afe_dat_1_0_filtered,
    output wire [13:0] afe_dat_1_1_filtered,
    output wire [13:0] afe_dat_1_2_filtered,
    output wire [13:0] afe_dat_1_3_filtered,
    output wire [13:0] afe_dat_1_4_filtered,
    output wire [13:0] afe_dat_1_5_filtered,
    output wire [13:0] afe_dat_1_6_filtered,
    output wire [13:0] afe_dat_1_7_filtered,
    output wire [13:0] afe_dat_1_8_filtered,
    output wire [13:0] afe_dat_2_0_filtered,
    output wire [13:0] afe_dat_2_1_filtered,
    output wire [13:0] afe_dat_2_2_filtered,
    output wire [13:0] afe_dat_2_3_filtered,
    output wire [13:0] afe_dat_2_4_filtered,
    output wire [13:0] afe_dat_2_5_filtered,
    output wire [13:0] afe_dat_2_6_filtered,
    output wire [13:0] afe_dat_2_7_filtered,
    output wire [13:0] afe_dat_2_8_filtered,
    output wire [13:0] afe_dat_3_0_filtered,
    output wire [13:0] afe_dat_3_1_filtered,
    output wire [13:0] afe_dat_3_2_filtered,
    output wire [13:0] afe_dat_3_3_filtered,
    output wire [13:0] afe_dat_3_4_filtered,
    output wire [13:0] afe_dat_3_5_filtered,
    output wire [13:0] afe_dat_3_6_filtered,
    output wire [13:0] afe_dat_3_7_filtered,
    output wire [13:0] afe_dat_3_8_filtered,
    output wire [13:0] afe_dat_4_0_filtered,
    output wire [13:0] afe_dat_4_1_filtered,
    output wire [13:0] afe_dat_4_2_filtered,
    output wire [13:0] afe_dat_4_3_filtered,
    output wire [13:0] afe_dat_4_4_filtered,
    output wire [13:0] afe_dat_4_5_filtered,
    output wire [13:0] afe_dat_4_6_filtered,
    output wire [13:0] afe_dat_4_7_filtered,
    output wire [13:0] afe_dat_4_8_filtered,
    input wire oeiclk,
    input wire fclk,
    output wire [31:0] dout,
    output wire [3:0] kout,
    input wire [31:0] Rcount_addr,
    output wire [63:0] Rcount
);

    st40_top st_wrapper(
        .reset_aclk(reset_aclk),
        .reset_fclk(reset_fclk),
        .adhoc(adhoc),
        .st_config(st_config),
        .signal_delay(signal_delay),
        .threshold_xc(threshold_xc),
        .ti_trigger(ti_trigger),
        .ti_trigger_stbr(ti_trigger_stbr),
        .reset_st_counters(reset_st_counters),
        .slot_id(slot_id),
        .crate_id(crate_id),
        .detector_id(detector_id),
        .version_id(version_id),
        .enable(enable),
        .afe_comp_enable(afe_comp_enable),
        .invert_enable(invert_enable),
        .st_40_signals_enable_reg(st_40_signals_enable_reg),
        .st_40_selftrigger_4_spybuffer(st_40_selftrigger_4_spybuffer),
        .filter_output_selector(filter_output_selector),
        .aclk(aclk),
        .timestamp(timestamp),
        .afe_dat_0_0(afe_dat_0_0),
        .afe_dat_0_1(afe_dat_0_1),
        .afe_dat_0_2(afe_dat_0_2),
        .afe_dat_0_3(afe_dat_0_3),
        .afe_dat_0_4(afe_dat_0_4),
        .afe_dat_0_5(afe_dat_0_5),
        .afe_dat_0_6(afe_dat_0_6),
        .afe_dat_0_7(afe_dat_0_7),
        .afe_dat_0_8(afe_dat_0_8),
        .afe_dat_1_0(afe_dat_1_0),
        .afe_dat_1_1(afe_dat_1_1),
        .afe_dat_1_2(afe_dat_1_2),
        .afe_dat_1_3(afe_dat_1_3),
        .afe_dat_1_4(afe_dat_1_4),
        .afe_dat_1_5(afe_dat_1_5),
        .afe_dat_1_6(afe_dat_1_6),
        .afe_dat_1_7(afe_dat_1_7),
        .afe_dat_1_8(afe_dat_1_8),
        .afe_dat_2_0(afe_dat_2_0),
        .afe_dat_2_1(afe_dat_2_1),
        .afe_dat_2_2(afe_dat_2_2),
        .afe_dat_2_3(afe_dat_2_3),
        .afe_dat_2_4(afe_dat_2_4),
        .afe_dat_2_5(afe_dat_2_5),
        .afe_dat_2_6(afe_dat_2_6),
        .afe_dat_2_7(afe_dat_2_7),
        .afe_dat_2_8(afe_dat_2_8),
        .afe_dat_3_0(afe_dat_3_0),
        .afe_dat_3_1(afe_dat_3_1),
        .afe_dat_3_2(afe_dat_3_2),
        .afe_dat_3_3(afe_dat_3_3),
        .afe_dat_3_4(afe_dat_3_4),
        .afe_dat_3_5(afe_dat_3_5),
        .afe_dat_3_6(afe_dat_3_6),
        .afe_dat_3_7(afe_dat_3_7),
        .afe_dat_3_8(afe_dat_3_8),
        .afe_dat_4_0(afe_dat_4_0),
        .afe_dat_4_1(afe_dat_4_1),
        .afe_dat_4_2(afe_dat_4_2),
        .afe_dat_4_3(afe_dat_4_3),
        .afe_dat_4_4(afe_dat_4_4),
        .afe_dat_4_5(afe_dat_4_5),
        .afe_dat_4_6(afe_dat_4_6),
        .afe_dat_4_7(afe_dat_4_7),
        .afe_dat_4_8(afe_dat_4_8),
        .afe_dat_0_0_filtered(afe_dat_0_0_filtered),
        .afe_dat_0_1_filtered(afe_dat_0_1_filtered),
        .afe_dat_0_2_filtered(afe_dat_0_2_filtered),
        .afe_dat_0_3_filtered(afe_dat_0_3_filtered),
        .afe_dat_0_4_filtered(afe_dat_0_4_filtered),
        .afe_dat_0_5_filtered(afe_dat_0_5_filtered),
        .afe_dat_0_6_filtered(afe_dat_0_6_filtered),
        .afe_dat_0_7_filtered(afe_dat_0_7_filtered),
        .afe_dat_0_8_filtered(afe_dat_0_8_filtered),
        .afe_dat_1_0_filtered(afe_dat_1_0_filtered),
        .afe_dat_1_1_filtered(afe_dat_1_1_filtered),
        .afe_dat_1_2_filtered(afe_dat_1_2_filtered),
        .afe_dat_1_3_filtered(afe_dat_1_3_filtered),
        .afe_dat_1_4_filtered(afe_dat_1_4_filtered),
        .afe_dat_1_5_filtered(afe_dat_1_5_filtered),
        .afe_dat_1_6_filtered(afe_dat_1_6_filtered),
        .afe_dat_1_7_filtered(afe_dat_1_7_filtered),
        .afe_dat_1_8_filtered(afe_dat_1_8_filtered),
        .afe_dat_2_0_filtered(afe_dat_2_0_filtered),
        .afe_dat_2_1_filtered(afe_dat_2_1_filtered),
        .afe_dat_2_2_filtered(afe_dat_2_2_filtered),
        .afe_dat_2_3_filtered(afe_dat_2_3_filtered),
        .afe_dat_2_4_filtered(afe_dat_2_4_filtered),
        .afe_dat_2_5_filtered(afe_dat_2_5_filtered),
        .afe_dat_2_6_filtered(afe_dat_2_6_filtered),
        .afe_dat_2_7_filtered(afe_dat_2_7_filtered),
        .afe_dat_2_8_filtered(afe_dat_2_8_filtered),
        .afe_dat_3_0_filtered(afe_dat_3_0_filtered),
        .afe_dat_3_1_filtered(afe_dat_3_1_filtered),
        .afe_dat_3_2_filtered(afe_dat_3_2_filtered),
        .afe_dat_3_3_filtered(afe_dat_3_3_filtered),
        .afe_dat_3_4_filtered(afe_dat_3_4_filtered),
        .afe_dat_3_5_filtered(afe_dat_3_5_filtered),
        .afe_dat_3_6_filtered(afe_dat_3_6_filtered),
        .afe_dat_3_7_filtered(afe_dat_3_7_filtered),
        .afe_dat_3_8_filtered(afe_dat_3_8_filtered),
        .afe_dat_4_0_filtered(afe_dat_4_0_filtered),
        .afe_dat_4_1_filtered(afe_dat_4_1_filtered),
        .afe_dat_4_2_filtered(afe_dat_4_2_filtered),
        .afe_dat_4_3_filtered(afe_dat_4_3_filtered),
        .afe_dat_4_4_filtered(afe_dat_4_4_filtered),
        .afe_dat_4_5_filtered(afe_dat_4_5_filtered),
        .afe_dat_4_6_filtered(afe_dat_4_6_filtered),
        .afe_dat_4_7_filtered(afe_dat_4_7_filtered),
        .afe_dat_4_8_filtered(afe_dat_4_8_filtered),
        .oeiclk(oeiclk),
        .fclk(fclk),
        .dout(dout),
        .kout(kout),
        .Rcount_addr(Rcount_addr),
        .Rcount(Rcount)
    );
endmodule